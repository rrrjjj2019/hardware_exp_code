`timescale 1ns/1ps

module Comparator_3bits (a, b, a_lt_b, a_gt_b, a_eq_b);
input [3-1:0] a, b;
output a_lt_b, a_gt_b, a_eq_b;

endmodule
