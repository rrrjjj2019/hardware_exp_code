`timescale 1ns/1ps

module Mux_8bits (a, b, sel, f);
input [8-1:0] a, b;
input sel;
output [8-1:0] f;

endmodule
