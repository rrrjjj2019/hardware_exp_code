    Mac OS X            	   2   �                                           ATTR         �   L                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine �[�[    �W    q/0083;5bfc4cf3;Safari;F8109516-6890-44DF-AD95-806784A17286 